//Name: EdgeDetector.sv
//Date: 2/13/2017
//Author: Omkar Pradhan
//Derived from: Dave Sluitter's 'majority.sv' module
//Description: This module detects positive and negative edge at the input (D) and outputs
// a short pulse at the ouput (posEdge and negEdge for positive edge and negative edge at D respectively)
